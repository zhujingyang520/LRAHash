// =============================================================================
// Module name: MemAccess
//
// This module exports the memory access stage of the computation datapath.
// =============================================================================

`include "pe.vh"

module MemAccess (
  input wire                  clk,              // system clock
  input wire                  rst,              // system reset

  // Input datapath & control path (memory stage)
  input wire                  comp_en_mem,      // computation enable (mem)
  input wire  [`PeDataBus]    in_act_value_mem, // input activation value (mem)
  input wire  [`PeActNoBus]   out_act_addr_mem, // output activation address
  input wire                  w_mem_cen,        // weight memory enable
  input wire                  w_mem_wen,        // weight memory write enable
  input wire  [`WMemAddrBus]  w_mem_addr,       // weight memory address

  // Output datapath & control path (mult stage)
  output reg                  comp_en_mult,     // computation enable (mult)
  output reg  [`PeDataBus]    in_act_value_mult,// input activation value (mult)
  output reg  [`PeDataBus]    w_value_mult,     // weight value (mult)
  output reg  [`PeActNoBus]   out_act_addr_mult // output activation address
);

// ---------------------
// Memory data output
// ---------------------
wire [`PeDataBus] w_mem_q;

// ----------------------------------------------------------------
// Instantiate the on-chip SRAM
// Note: The memory model is generated by CACTI 6.5
// - W Memory size: 16x65536
// ----------------------------------------------------------------
`ifdef CACTI_MEM_MODEL
// memory output enable (active low)
reg w_mem_oe;
always @ (posedge clk or posedge rst) begin
  if (rst) begin
    w_mem_oe          <= 1'b1;
  end else begin
    w_mem_oe          <= w_mem_cen;
  end
end
// memory behavior model generated by `cacti-mc`
SRAM_16x65536_1P w_mem (
  .CE1                (clk),                    // system clock
  .WEB1               (w_mem_wen),              // write enable (active low)
  .CSB1               (w_mem_cen),              // chip enable (active low)
  .OEB1               (w_mem_oe),               // output enable (active low)
  .A1                 (w_mem_addr),             // read/write address
  .I1                 (`W_MEM_ADDR_WIDTH'd0),   // data input (write op)
  .O1                 (w_mem_q)                 // data output (read op)
);
`else
// ideal memory model (WARNING: not synthesizable!)
spram_behav # (
  .MEM_WIDTH          (`W_MEM_DATA_WIDTH),      // memory (bus) width
  .MEM_DEPTH          (2**`W_MEM_ADDR_WIDTH)    // memory depth
) w_mem (
  .clk                (clk),                    // system clock
  .cen                (w_mem_cen),              // chip enable (active low)
  .wen                (w_mem_wen),              // write enable (active low)
  .addr               (w_mem_addr),             // read/write address
  .d                  (`W_MEM_ADDR_WIDTH'd0),   // data input (write op)
  .q                  (w_mem_q)                 // data output (read op)
);
`endif

// ----------------------------------------------
// Pipeline stage of the datapath & control path
// ----------------------------------------------
always @ (posedge clk or posedge rst) begin
  if (rst) begin
    comp_en_mult      <= 1'b0;
    in_act_value_mult <= 0;
    out_act_addr_mult <= 0;
    w_value_mult      <= 0;
  end else begin
    comp_en_mult      <= comp_en_mem;
    in_act_value_mult <= in_act_value_mem;
    out_act_addr_mult <= out_act_addr_mem;
    w_value_mult      <= w_mem_q;
  end
end

endmodule
